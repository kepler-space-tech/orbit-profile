--------------------------------------------------------------------------------
-- Project: {{ orbit.ip }}
-- Author:  {{ orbit.user }}
-- Entity:  {{ orbit.ip.name }}
-- Created: {{ orbit.date }}
-- Details:
--
--
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity {{ orbit.ip.name }} is
    generic(

    );
    port(

    );
end entity {{ orbit.ip.name }};


architecture rtl of {{ orbit.ip.name }} is

begin


end architecture rtl;