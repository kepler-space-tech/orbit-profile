--------------------------------------------------------------------------------
-- Project: {{ orbit.ip }}
-- Author:  {{ orbit.user }}
-- Entity:  {{ orbit.filename}}
-- Created: {{ orbit.date }}
-- Details:
--
--
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity {{ orbit.filename }} is
    generic(

    );
    port(

    );
end entity {{ orbit.filename }};


architecture rtl of {{ orbit.filename }} is

begin


end architecture rtl;